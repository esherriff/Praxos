library ieee;
use ieee.std_logic_1164.all;

-- Praxos ROM content

package praxos_application_image is

	type application_image_t is array(0 to (2**8)-1) of std_logic_vector(35 downto 0);
	constant application_image : application_image_t := (
		0 =>"001100000000000000000000000000000001", -- 0 			LD#	1
		1 =>"011000000000000000000000000000000001", -- 1 			ST	SCRATCH
		2 =>"001000000000000000000000000000000000", -- 2 			ILD#	0
		3 =>"001100000000000000000000000000001010", -- 3 @MAIN	LD#	DEC
		4 =>"101100001111111111111111111111111111", -- 4 			JAL	CALL
		5 =>"010000000000000000000000000000000010", -- 5 			LD	IO
		6 =>"010011000000000000000000000000000001", -- 6 			XOR	SCRATCH
		7 =>"011000000000000000000000000000000010", -- 7 			ST	IO
		8 =>"010100000000000000000000000000000000", -- 8 			OUT	0
		9 =>"111000011111111111111111111111111001", -- 9 			BRA	MAIN
		10 =>"110100000000000000000000000000000000", -- 10 @DEC		DECI
		11 =>"001100000000000000000000000000000101", -- 11 			LD#	5
		12 =>"000010100000000000000000000000000001", -- 12 @DEC_LP	SUB#	1
		13 =>"111001011111111111111111111111111110", -- 13 			BRNZ	DEC_LP
		14 =>"110000000000000000000000000000000000", -- 14 			LDI	0
		15 =>"100100000000000000000000000000000000", -- 15 			INCI
		16 =>"101100001111111111111111111111111111", -- 16 			JAL	RET
		17 =>"111011100000000000000000000000000000", -- 17 			NOP
		others => (others => '0'));
end praxos_application_image;
